-- State machine