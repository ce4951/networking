-- Timer